
 
interface mux_if;
 logic [3:0] a;
 logic [3:0] b;
 logic [3:0] c;
 logic [3:0] d;
 logic [1:0] sel;
 logic [3:0] y;
endinterface
