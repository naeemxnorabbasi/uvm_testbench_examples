////////////////////////////////////////////////////////////
 
interface spi_i;
 
   logic clk, rst, cs, miso;
   logic ready, mosi, op_done;
    
endinterface
