
interface add_if;
 logic [3:0] add_in1,add_in2;
 logic clk, rst;
 logic [4:0] add_out;
endinterface
 
 
//////////////////////////////
 
interface mul_if;
 logic [3:0] mul_in1,mul_in2;
 logic clk, rst;
 logic [7:0] mul_out;
endinterface
 
////////////////////////////////////////
 
