package pipe_pkg;

   import uvm_pkg::*;

`include "uvm_macros.svh"
`include "data_packet.sv"
`include "driver.sv"
`include "monitor.sv"
`include "sequencer.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "pipe_coverage.sv"
`include "pipe_env.sv"
`include "dut_env.sv"
`include "pipe_sequence_lib.sv"
`include "test_lib.sv"   
   
endpackage // pipe_pkg
   
